library ieee;
use ieee.std_logic_1164.all;

entity myAnd is
  
  port (
    myBtn_1 : in  std_logic;
    myBtn_2 : in  std_logic;
    myOut   : out std_logic);

end entity myAnd;
