architecture rtl of myAnd is

begin

  myOut <= (not myBtn_1) and (not myBtn_2);

end architecture rtl;

